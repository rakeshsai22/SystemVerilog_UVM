package jtag_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"
`include "jtag_interface.sv"
`include "jtag_seq_item.sv"
`include "jtag_sqr.sv"
`include "jtag_drv.sv"
`include "jtag_mon.sv"
`include "jtag_agent.sv"
`include "jtag_env.sv"
`include "jtag_seq.sv"
`include "jtag_test.sv"
// `include "jtag_packet.sv"


endpackage