// functions test

// testbench