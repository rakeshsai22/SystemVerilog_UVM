// write a constraint to generate two consecutive 1's in a 16 bit variable

class pkt;
  rand bit [15:0] a;
  constraint c
