interface fulladd_if(input logic clk);
  logic [3:0] a ;
  logic [3:0] b ;
  logic c_in ;
  reg c_out ;
  reg [3:0] sum ;
endinterface