interface synchronous_counter_if(input logic clk);
  logic rst_n ;
  logic up ;
  logic [SIZE-1:0] cnt ;
endinterface