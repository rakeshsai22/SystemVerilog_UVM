// to generate unique values for the variables/elements in an array (fixed array, associative array, dynamic array, queue, stack, list, etc)

// syntax : constraint <name> {unique {array or varuiable name};}

typedef enum  { r,a,n,d,o,m } scale_e;

class seq_item;
    rand bit [3:0] arr_s[5];
    rand bit [3:0] arr_d[];
    rand
    
endclass