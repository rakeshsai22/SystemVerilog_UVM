interface jtag_if;
  logic TCK;
  logic TDI;
  logic TMS;
  logic TRST_N;
  logic TDO;
endinterface
