module fifo_syn #(
    parameter FIFO_DEPTH = 8;
    parameter DATA_WIDTH = 32
) (
    
);
    
endmodule