package fulladd_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "fulladd_seq_item.sv"
  `include "fulladd_seq.sv"
  `include "fulladd_sequencer.sv"
  `include "fulladd_driver.sv"
  `include "fulladd_monitor.sv"
  `include "fulladd_agent.sv"
  `include "fulladd_env.sv"
  `include "fulladd_test.sv"

endpackage : fulladd_pkg