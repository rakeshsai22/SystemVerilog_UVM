// functions test

