// mailbox is a way to allow different processes to exchange data betwen each other
//  created with a bounded or unbounded queue size
// ## teo types of mailboxes 
//      1. Generic - accepts any data type
