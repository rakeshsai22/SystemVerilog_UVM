// Virtual methods

// a virtual method or task from the base class can be overridden by a method of its child class having the same method name and arguments

// ?? virtual class / abstract class 



