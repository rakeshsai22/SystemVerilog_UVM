// Associative array stores entries in a sparse matrix format. 
// these arrs allocate the storage only when it is used, unless like in the dynamic array where the storage is allocated at the time of declaration.
// the index expression is not restricted to a simple integer or string, it can be any data type.
// Associative arrays are not allowed in the class, they can be declared only in the module or program block.
// Associative array implements a lookup table of the elements of its declared type. The data type to be used as an index serves as lookup key and imposes an ordering

//  Usage : When the size of the collection is unknown or the data space is sparse.

// data_type array_name [index_type] ;